
/****************************************************************************
 * SVParamVal.svh
 ****************************************************************************/

  
/**
 * Class: SVParamVal
 * 
 * TODO: Add class documentation
 */
class SVParamVal extends IParamVal ;

	function new();

	endfunction


endclass


