
/****************************************************************************
 * IInterfaceInst.svh
 ****************************************************************************/

  
/**
 * Class: IInterfaceInst
 * 
 * TODO: Add class documentation
 */
class IInterfaceInst;
	chandle			m_hndl;
		
endclass


