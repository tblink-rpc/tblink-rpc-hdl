
/****************************************************************************
 * DpiTbLinkListener.svh
 ****************************************************************************/

  
/**
 * Class: DpiTbLinkListener
 * 
 * TODO: Add class documentation
 */
class DpiTbLinkListener;

	function new();

	endfunction


endclass


