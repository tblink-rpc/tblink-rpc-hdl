/****************************************************************************
 * IParamValStr.svh
 ****************************************************************************/

  
/**
 * Class: IParamValStr
 * 
 * TODO: Add class documentation
 */
class IParamValStr extends IParamVal;

	virtual function string val();
		return "";
	endfunction

endclass


