
/****************************************************************************
 * IInterfaceType.svh
 ****************************************************************************/

  
/**
 * Class: IInterfaceType
 * 
 * TODO: Add class documentation
 */
class IInterfaceType;
	
endclass

