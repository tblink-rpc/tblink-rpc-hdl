
/****************************************************************************
 * IInterfaceType.svh
 ****************************************************************************/

  
/**
 * Class: IInterfaceType
 * 
 * TODO: Add class documentation
 */
class IInterfaceType;
	chandle			m_hndl;
endclass

