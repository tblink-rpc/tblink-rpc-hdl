/****************************************************************************
 * DpiTypeMap.svh
 ****************************************************************************/

  
/**
 * Class: DpiTypeMap
 * 
 * TODO: Add class documentation
 */
class DpiTypeMap extends ITypeMap;
	chandle			m_hndl;

	function new(chandle hndl);
		m_hndl = hndl;
	endfunction

endclass


