/****************************************************************************
 * SvInterfaceTypeBuilder.svh
 ****************************************************************************/

  
/**
 * Class: SvInterfaceTypeBuilder
 * 
 * TODO: Add class documentation
 */
class SvInterfaceTypeBuilder extends IInterfaceTypeBuilder;

	function new();

	endfunction


endclass


