
/****************************************************************************
 * IParamValInt.svh
 ****************************************************************************/

  
/**
 * Class: IParamValInt
 * 
 * TODO: Add class documentation
 */
class IParamValInt extends IParamVal;
		
endclass

