/****************************************************************************
 * ITypeVec.svh
 ****************************************************************************/

  
/**
 * Class: ITypeVec
 * 
 * TODO: Add class documentation
 */
class ITypeVec extends IType;

	virtual function IType elem_t();
		return null;
	endfunction

endclass


