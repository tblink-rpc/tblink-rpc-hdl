
/****************************************************************************
 * IParamValMap.svh
 ****************************************************************************/

  
/**
 * Class: IParamValMap
 * 
 * TODO: Add class documentation
 */
class IParamValMap extends IParamVal;
endclass


