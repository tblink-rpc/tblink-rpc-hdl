
/****************************************************************************
 * DpiInterfaceType.svh
 ****************************************************************************/

  
/**
 * Class: DpiInterfaceType
 * 
 * TODO: Add class documentation
 */
class DpiInterfaceType extends IInterfaceType;
	chandle				m_hndl;

	function new(chandle hndl);
		m_hndl = hndl;
	endfunction


endclass


