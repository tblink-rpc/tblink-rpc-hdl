
/****************************************************************************
 * IMethodTypeBuilder.svh
 ****************************************************************************/

  
/**
 * Class: IMethodTypeBuilder
 * 
 * TODO: Add class documentation
 */
class IMethodTypeBuilder;

	virtual function void add_param(
		string					name,
		IType					ptype);
	endfunction

endclass


