
/****************************************************************************
 * SVInvokeInfo.svh
 ****************************************************************************/

  
/**
 * Class: SVInvokeInfo
 * 
 * TODO: Add class documentation
 */
class SVInvokeInfo extends InvokeInfo;

	function new();

	endfunction


endclass


