/****************************************************************************
 * tblink_rpc_uvm.sv
 ****************************************************************************/
`include "uvm_macros.svh"
  
/**
 * Package: tblink_rpc_uvm
 * 
 * TODO: Add package documentation
 */
package tblink_rpc_uvm;
	import uvm_pkg::*;
	import tblink_rpc::*;


endpackage


