
/****************************************************************************
 * IParamValInt.svh
 ****************************************************************************/

  
/**
 * Class: IParamValInt
 * 
 * TODO: Add class documentation
 */
class IParamValInt extends IParamVal;
	
	virtual function longint val_s();
	endfunction
	
	virtual function longint unsigned val_u();
	endfunction
		
endclass

