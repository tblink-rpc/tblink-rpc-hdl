
/****************************************************************************
 * IParamValBool.svh
 ****************************************************************************/

  
/**
 * Class: IParamValBool
 * 
 * TODO: Add class documentation
 */
class IParamValBool extends IParamVal;
		
	virtual function bit val();
		return 0;
	endfunction
		
endclass


