/****************************************************************************
 * tblink_rpc_uvm.sv
 ****************************************************************************/
`include "uvm_macros.svh"
  
/**
 * Package: tblink_rpc_uvm
 * 
 * TODO: Add package documentation
 */
package tblink_rpc_uvm;
	import uvm_pkg::*;
	import tblink_rpc::*;

	`include "TbLinkAgentConfig.svh"
	`include "TbLinkAgent.svh"
	`include "TbLinkLaunchSeqBase.svh"
	`include "TbLinkLaunchSeq.svh"
	
	`include "TbLinkLaunchUvmObj.svh"
	`include "TbLinkLaunchUvmSeq.svh"


endpackage


