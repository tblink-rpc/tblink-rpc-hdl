/****************************************************************************
 * uvm_python_pkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"
  
/**
 * Package: uvm_python_pkg
 * 
 * TODO: Add package documentation
 */
package uvm_python_pkg;
	import uvm_pkg::*;
	import tblink_rpc::*;
	import tblink_rpc_uvm::*;

	`include "uvm_python_seq_if.svh"
	`include "uvm_python_remote_obj.svh"
	
	`include "uvm_python_test.svh"


endpackage


