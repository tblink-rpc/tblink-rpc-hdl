
/****************************************************************************
 * DpiTypeVec.svh
 ****************************************************************************/

  
/**
 * Class: DpiTypeVec
 * 
 * TODO: Add class documentation
 */
class DpiTypeVec extends ITypeVec;
	chandle			m_hndl;

	function new(chandle hndl);
		m_hndl = hndl;
	endfunction

endclass


